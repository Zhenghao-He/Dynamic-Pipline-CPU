`define COND_FLOW 2'b00
`define COND_STALL 2'b01
`define COND_ZERO 2'b10
`define PC_ADDR_INIT 32'h00400000
`define IR_NON 32'hffffffff
`define IR_NON_31_26 6'b111111
`define MULU 2'b00
`define MUL 2'b01
`define DIVU 2'b10
`define DIV 2'b11
`define EXTEND5_Z 3'b000
`define EXTEND16_SL2_S 3'b001
`define EXTEND16_Z 3'b010
`define EXTEND16_S 3'b011
`define EXTEND8_Z 3'b100
`define EXTEND8_S 3'b101
`define EXTEND32_NON 3'b110
`define SELECT_PC_NPCEXT 3'b000
`define SELECT_PC_RS 3'b001
`define SELECT_PC_INTR_ADDR 3'b010
`define SELECT_PC_EPC 3'b011
`define SELECT_PC_CONNECT 3'b100
`define SELECT_PC_NPC 3'b101
`define SELECT_ALUa_HI 3'b000
`define SELECT_ALUa_LO 3'b001
`define SELECT_ALUa_NPC 3'b010
`define SELECT_ALUa_RS 3'b011
`define SELECT_ALUa_EXT 3'b100
`define SELECT_ALUa_CP0 3'b101
`define SELECT_ALUa_IMM0 3'b110
`define SELECT_ALUb_IMM0 2'b00
`define SELECT_ALUb_RT 2'b01
`define SELECT_ALUb_EXT 2'b10
`define SELECT_RDC_IR_15_11 2'b00
`define SELECT_RDC_IR_20_16 2'b01
`define SELECT_RDC_IMM31 2'b10
`define SELECT_RD_Z 2'b00
`define SELECT_RD_MEM 2'b01
`define SELECT_RD_HI 2'b10
`define SELECT_RD_LO 2'b11
`define WIDTH_32 2'b00
`define WIDTH_16 2'b01
`define WIDTH_8 2'b10
`define NORMAL 2'b00
`define OVERFLOW 2'b01
`define MULDIV 2'b10
`define VIOLATE 2'b11

